module data_mem(
	input wire clk,
	input wire mem_read,
	input wire mem_write,
	input wire 
